module led_output(
	input clk,
	input [7:0] data,
	output [7:0] LED);
	
	
	always@(c
	
endmodule