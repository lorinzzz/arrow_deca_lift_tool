// selects between the active_buzzer_light_sensor or the active_buzzer_gsensor circuit

module buzzer_multiplxer()